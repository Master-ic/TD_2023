module speed_up( );



endmodule
